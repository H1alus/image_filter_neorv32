-- ================================================================================ --
-- image_filter_NEORV32: hardware accelerated image filter for neorv32              --                
-- -------------------------------------------------------------------------------- --
-- Project repository - https://github.com/H1alus/image_filter_neorv32              --
-- Copyright (c) 2024 Vittorio Folino. All rights reserved.                         --
-- Licensed under the BSD-3-Clause license, see LICENSE for details.                --
-- SPDX-License-Identifier: BSD-3-Clause                                            --
-- ================================================================================ --
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

library std;
use std.textio.all;
use std.env.finish;

library neorv32;
use neorv32.neorv32_package.all;
use neorv32.neorv32_application_image.all; -- this file is generated by the image generator

entity neorv32_tb is
--  Port ( );
end neorv32_tb;

architecture Behavioral of neorv32_tb is
  constant f_clock_c               : natural := 100_000_000; --clock frequency of the uut
  constant baud0_rate_c            : natural := 19200; -- simulation UART0 (primary UART) baud rate
  -- internals - hands off! --
  constant uart0_baud_val_c : real := real(f_clock_c) / real(baud0_rate_c);
  constant t_clock_c        : time := (1 sec) / f_clock_c;
  -- generators --
  signal clk_gen, rstn_gen : std_ulogic := '0';
  -- uart --
  signal uart0_txd : std_ulogic;
  
  -- maximum memory size in bytes --
  constant MEM_SIZE : natural := 8*1024; -- total memory size in bytes
  constant MEM_FILE : string := "/mnt/shared/inputfile.txt";
  
  -- [NOTE] sizes >= 4MB are crashing GHDL in this setup; maximum still-OK-size = 3MB
  constant mem_size_max_c : natural := 2*1024*1024; -- just use 2MB as maximum to be safe ;)

  -- make sure actual memory size is a power of two (or <mem_size_max_c> for the rare case or very large images) --
  constant mem_size_c : natural := cond_sel_natural_f(boolean(MEM_SIZE >= mem_size_max_c), mem_size_max_c, 2**index_size_f(MEM_SIZE));
  
  -- memory type --
  type mem8_bv_t is array (natural range <>) of std_logic_vector(7 downto 0); -- bit_vector type for optimized system storage
  
  -- initialize mem8_bv_t array from plain ASCII HEX file  --
  impure function mem8_bv_init_f(file_name : string; num_bytes : natural; byte_sel : natural) return mem8_bv_t is
    file     text_file   : text open read_mode is file_name;
    variable text_line_v : line;
    variable mem8_bv_v   : mem8_bv_t(0 to num_bytes-1);
    variable index_v     : natural;
    variable word_v      : std_logic_vector(31 downto 0);
  begin
    mem8_bv_v := (others => (others => '0')); -- initialize to all-zero
    index_v   := 0;
    while (endfile(text_file) = false) and (index_v < num_bytes) loop
      readline(text_file, text_line_v);
      hread(text_line_v, word_v);
      case byte_sel is
        when 0      => mem8_bv_v(index_v) := word_v(07 downto 00);
        when 1      => mem8_bv_v(index_v) := word_v(15 downto 08);
        when 2      => mem8_bv_v(index_v) := word_v(23 downto 16);
        when others => mem8_bv_v(index_v) := word_v(31 downto 24);
      end case;
      index_v := index_v + 1;
    end loop;
    return mem8_bv_v;
  end function mem8_bv_init_f;


  -- memory address --
  signal addr : integer range 0 to (mem_size_c/4)-1;
  
  
  -- simulated external Wishbone memory C (can be used to simulate external IO access) --
  constant ext_mem_c_base_addr_c   : std_ulogic_vector(31 downto 0) := x"F0000000"; -- wishbone memory base address (default begin of EXTERNAL IO area)
  --constant ext_mem_c_size_c        : natural := 64*1024; -- wishbone memory size in bytes, should be smaller than an iCACHE block
  constant ext_mem_c_end_addr_c    : std_ulogic_vector(31 downto 0) := 
  std_ulogic_vector(to_unsigned(to_integer(unsigned(ext_mem_c_base_addr_c)) + mem_size_c, 32));
  
   -- Wishbone bus --
  type wishbone_t is record
    addr  : std_ulogic_vector(31 downto 0); -- address
    wdata : std_ulogic_vector(31 downto 0); -- master write data
    rdata : std_ulogic_vector(31 downto 0); -- master read data
    tag   : std_ulogic_vector(2 downto 0); -- access tag
    we    : std_ulogic; -- write enable
    sel   : std_ulogic_vector(3 downto 0); -- byte enable
    stb   : std_ulogic; -- strobe
    cyc   : std_ulogic; -- valid cycle
    ack   : std_ulogic; -- transfer acknowledge
    err   : std_ulogic; -- transfer error
  end record;
  signal wb_cpu : wishbone_t;
  signal first_ack : std_logic;
  
    -- Wishbone access latency type --
  type ext_mem_read_latency_t is array (0 to 255) of std_ulogic_vector(31 downto 0);

component neorv32_mine is
  port (
    -- Global control --
    clk_i  : in  std_logic;
    rstn_i : in  std_logic;
    
    -- External bus interface (available if XBUS_EN = true) --
    xbus_adr_o     : out std_ulogic_vector(31 downto 0);                    -- address
    xbus_dat_o     : out std_ulogic_vector(31 downto 0);                    -- write data
    xbus_tag_o     : out std_ulogic_vector(2 downto 0);                     -- access tag
    xbus_we_o      : out std_ulogic;                                        -- read/write
    xbus_sel_o     : out std_ulogic_vector(3 downto 0);                     -- byte enable
    xbus_stb_o     : out std_ulogic;                                        -- strobe
    xbus_cyc_o     : out std_ulogic;                                        -- valid cycle
    xbus_dat_i     : in  std_ulogic_vector(31 downto 0) := (others => 'L'); -- read data
    xbus_ack_i     : in  std_ulogic := 'L';                                 -- transfer acknowledge
    xbus_err_i     : in  std_ulogic := 'L';                                 -- transfer error
    
    -- primary UART0 (available if IO_UART0_EN = true) --
    uart0_txd_o    : out std_ulogic;                                        -- UART0 send data
    uart0_rxd_i    : in  std_ulogic;                                 -- UART0 receive data
    uart0_rts_o    : out std_ulogic;                                        -- HW flow control: UART0.RX ready to receive ("RTR"), low-active, optional
    uart0_cts_i    : in  std_ulogic;                                 -- HW flow control: UART0.TX allowed to transmit, low-active, optional

--    -- CPU interrupts (for chip-internal usage only) --
    mtime_irq_i    : in  std_ulogic := 'L';                                 -- machine timer interrupt, available if IO_MTIME_EN = false
    msw_irq_i      : in  std_ulogic := 'L';                                 -- machine software interrupt
    mext_irq_i     : in  std_ulogic := 'L'                                  -- machine external interrupt
  );
end component;
  
  component uart_rx is
  generic (
    name : string;
    uart_baud_val_c : real);

    port (
      clk : in std_ulogic;
      uart_txd : in std_ulogic
     );
  end component;

  file file_uart_tx_out : text open write_mode is "neorv32.testbench_uart0.out";

begin

  
  -- Clock/Reset Generator ------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------

  clk_gen <= not clk_gen after (t_clock_c/2);
  rstn_gen <= '0', '1' after 200*(t_clock_c/2);
  
  -- The core of the problem -----------------------------------------------------------------
  -- -----------------------------------------------------------------------------------------
  uut: neorv32_mine
  port map(    
     -- Global control --
    clk_i  => clk_gen,    -- global clock, rising edge
    rstn_i => rstn_gen,   -- global reset, low-active, async
    -- PWM (available if IO_PWM_NUM_CH > 0) --
    
    -- primary UART0 (available if IO_UART0_EN = true) --
    uart0_txd_o    => uart0_txd,       -- UART0 send data
    uart0_rxd_i => uart0_txd,
    uart0_cts_i    => '0',       -- HW flow control: UART0.TX allowed to transmit, low-active, optional

     -- External bus interface (available if XBUS_EN = true) --
    xbus_adr_o     => wb_cpu.addr,     -- address
    xbus_dat_o     => wb_cpu.wdata,    -- write data
    xbus_tag_o     => wb_cpu.tag,      -- access tag
    xbus_we_o      => wb_cpu.we,       -- read/write
    xbus_sel_o     => wb_cpu.sel,      -- byte enable
    xbus_stb_o     => wb_cpu.stb,      -- strobe
    xbus_cyc_o     => wb_cpu.cyc,      -- valid cycle
    xbus_dat_i     => wb_cpu.rdata,    -- read data
    xbus_ack_i     => wb_cpu.ack,      -- transfer acknowledge
    xbus_err_i     => wb_cpu.err      -- transfer error
  );
  
 -- UART Simulation Receiver ---------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  uart0_checker: uart_rx
  generic map (
    name => "uart0",
    uart_baud_val_c => uart0_baud_val_c
  )
  port map (
    clk => clk_gen,
    uart_txd => uart0_txd
  );

  -- External Main Memory [rwx] - Constructed from four parallel byte-wide memories ---------
  -- -------------------------------------------------------------------------------------------
  ext_mem_rw: process(clk_gen)
    file outfile : text open write_mode is "/mnt/shared/ram_1.txt";
    variable lined_v : line;
    variable mem8_bv_b0_v : mem8_bv_t(0 to (mem_size_c/4)-1) := mem8_bv_init_f(MEM_FILE, mem_size_c/4, 0);
    variable mem8_bv_b1_v : mem8_bv_t(0 to (mem_size_c/4)-1) := mem8_bv_init_f(MEM_FILE, mem_size_c/4, 1);
    variable mem8_bv_b2_v : mem8_bv_t(0 to (mem_size_c/4)-1) := mem8_bv_init_f(MEM_FILE, mem_size_c/4, 2);
    variable mem8_bv_b3_v : mem8_bv_t(0 to (mem_size_c/4)-1) := mem8_bv_init_f(MEM_FILE, mem_size_c/4, 3);
  begin
    if rising_edge(clk_gen) then
       first_ack <= wb_cpu.stb;
       wb_cpu.ack <= first_ack and wb_cpu.cyc;
       wb_cpu.rdata <= (others => '0');
       wb_cpu.err <= '0';
      if first_ack and wb_cpu.cyc then
        if ( wb_cpu.we = '1') then -- byte-wide write access
          if ( wb_cpu.sel(0) = '1') then mem8_bv_b0_v(addr) := wb_cpu.wdata(07 downto 00); end if;
          if ( wb_cpu.sel(1) = '1') then mem8_bv_b1_v(addr) := wb_cpu.wdata(15 downto 08); end if;
          if ( wb_cpu.sel(2) = '1') then mem8_bv_b2_v(addr) := wb_cpu.wdata(23 downto 16); end if;
          if ( wb_cpu.sel(3) = '1') then mem8_bv_b3_v(addr) := wb_cpu.wdata(31 downto 24); end if;
          write(lined_v, "0x" & to_hstring(wb_cpu.wdata));
          writeline(outfile,lined_v);
          
        else -- word-aligned read access
          wb_cpu.rdata(07 downto 00) <= to_stdulogicvector(mem8_bv_b0_v(addr));
          wb_cpu.rdata(15 downto 08) <= to_stdulogicvector(mem8_bv_b1_v(addr));
          wb_cpu.rdata(23 downto 16) <= to_stdulogicvector(mem8_bv_b2_v(addr));
          wb_cpu.rdata(31 downto 24) <= to_stdulogicvector(mem8_bv_b3_v(addr));
        end if;
      end if;
    end if;
  end process ext_mem_rw;
  -- read/write address --

  addr <= to_integer(unsigned(wb_cpu.addr(index_size_f(mem_size_c/4)+1 downto 2)));

end Behavioral;
